*Summing Amplifier with Opamp 741 
*Opamp 741 contains 26 BJT
* Original freeda netlist by Muhammad Kabir
* Modifications: removed substrate connections (not used anyway) 
*                and dummy resistors

.options maxiter=100 gyr=1e-5 maxdelta=3. sparse=1
*.analysis op intvars=0
.analysis eop gcomp=.5mS 

xamp1 vplus vminus vout lm741
xmain1 vplus vminus vout extcircuit


# External circuit
.subckt extcircuit vplus vminus vout
vsin:v2 153 0 vdc=1. acmag=.1 rint = 5.
vpulse:v2 154 153 rint=5 v1=0 v2=2. pw=400us per=1ms td=50us tr=50us tf=50us
vsin:v1 151 0 mag=.2 freq=5kHz
res:r1s 151 152 r=10.

res:r1ext 152 vminus r=5e3
res:r2ext 154 vminus r=20e3
res:r4ext vminus 23 r=20e3
res:r5ext vplus 0 r=3.33e3
.ends


#####################################################################
.subckt lm741 201 202 23
*** OPAMP LM 741 ***

***Power Supply****
***VCC PIN 1
***VEE PIN 2

vdc:vcc 100 0 vdc=7.5
res:rcc 1 100 r=20
vdc:vee 0 101 vdc=7.5
res:ree 101 2 r=20

***Widlar Current Source***
svbjt:q10 5 4 3 model=mynpn area=1
svbjt:q11 4 4 2 model=mynpn area=1
res:r4 3 2 r=5e3
res:r5 6 4 r=39e3
svbjt:q9 5 7 1 model=mypnp area=1
svbjt:q12 6 6 1 model=mypnp area=1

svbjt:q13b 15 6 1 model=mypnp area=3
svbjt:q13a 16 6 1 model = mypnp area=1

svbjt:q8 7 7 1 model = mypnp area=1

***INPUT***
*Vplus ---> PIN201
*Vminus---> PIN202
*Offset null1 ----> PIN14
*Offset null2 ----> PIN17

***Differential Amplifier***
svbjt:q1 7 201 9 model = mynpn area=1
svbjt:q2 7 202 10 model = mynpn area=1
svbjt:q3 11 5 9 model = mypnp area=1
svbjt:q4 12 5 10 model = mypnp area=1
svbjt:q5 11 13 14 model = mynpn area=1
svbjt:q6 12 13 17 model = mynpn area=1
svbjt:q7 1 11 13 model = mynpn area=1
res:r1 14 2 r=1e3
res:r2 17 2 r=1e3
res:r3 13 2 r=50e3


svbjt:q19 16 16 20 model = mynpn area=1
svbjt:q18 16 20 21 model = mynpn area=1
res:r10 20 21 r=40e3
cap:cc 15 12 c=30e-12


svbjt:q16 1 12 18 model = mynpn area=1
svbjt:q17 15 18 19 model = mynpn area=1
svbjt:q22 12 25 2 model = mynpn area=1
res:r9 18 2 r=50e3
res:r8 19 2 r=100

svbjt:q23b 2 15 12 model = mypnp area=1
svbjt:q23a 2 15 21 model = mypnp area=1

***Output***
*Output ---> PIN23

svbjt:q14 1 16 22 model = mynpn area=3
svbjt:q15 16 22 23 model = mynpn area=1
res:r6 22 23 r=27
svbjt:q21 25 24 23 model = mypnp area=1
res:r7 23 24 r=22
svbjt:q20 2 21 24 area=1 type=pnp isat=1e-14 rb=150  \
br=4 bf=50 vaf=50 tf=20e-9 cje=0.5e-12 cjc=2e-12
* rc=50 re=2

svbjt:q24 25 25 2 model = mynpn area=1
res:r12 25 2 r=50e3

.model mynpn svbjt(type=npn isat=5e-15 rb=200 bf=200 \
br=2 vaf=130 tf=0.35e-9 cje=1e-12 cjc=0.3e-12 \
ne=0.33 nc=0.5 tr=400e-9 vje=0.7 vjc=0.55 rc=200 re=2)

.model mypnp svbjt(type=pnp isat=2e-15 rb=300 \
bf=50 br=4 vaf=50 tf=30e-9 cje=0.3e-12 cjc=1e-12 \
ne=0.5 nc=0.5 tr=3000e-9 vje=0.55 vjc=0.55 rc=100  re=10)

.ends
#####################################################################

.end
